library verilog;
use verilog.vl_types.all;
entity Processador_mips_final_vlg_vec_tst is
end Processador_mips_final_vlg_vec_tst;
