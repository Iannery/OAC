library verilog;
use verilog.vl_types.all;
entity memMIPS_vlg_vec_tst is
end memMIPS_vlg_vec_tst;
